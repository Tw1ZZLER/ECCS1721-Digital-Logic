-------------------------------------------------------------------------------------
-- Transceiver Hardware Component Container, version 2 (for Mk8 Apex/XCVR)
-------------------------------------------------------------------------------------
-- Author:      Maxwell Phillips
-- Copyright:   Ohio Northern University, 2023.
-- License:     GPL v3
-- Description: Container for hardware to be wrapped by apex component.
-------------------------------------------------------------------------------------
--
-- This file is the hardware component container wrapped by the top level apex
-- component. You should modify this file to wrap your hardware in order to utilize
-- it with the serial transceiver. See the apex component and transceiver files
-- for more details on their functionality.
--
-------------------------------------------------------------------------------------
-- Generics
-------------------------------------------------------------------------------------
--
-- [G_byte_bits]: Should be 8. Mapped from top-level component.
--
-- [G_total_bits]: The capacity, in bits, of the transceiver.
--                 Mapped directly from the top-level component.
--                 Should be used to help structure hardware components.
--
-- [G_clk_freq]: Should match the clock frequency of the FPGA board.
--               Again, mapped by top-level component.
--
-------------------------------------------------------------------------------------
-- Ports
-------------------------------------------------------------------------------------
--
-- [clk_100mhz]: Input clock signal; should match [G_clk_freq] generic.
--
-- [clk_hw]: Clock signal to time contained hardware. Generated by MMCM on top-level.
--
-- [reset]: Asynchronous reset signal. The module should be initially
--          reset automatically by the transceiver, and will remain reset
--          until all bytes are received and the processing stage begins.
--          To preserve state, the hardware is NOT reset after the processing
--          stage and during the transmission stage. This allows displaying
--          output on the LEDs from the hardware container more easily.
--
-- [load]: Signal which is received for one clock cycle (of [G_clk_freq]) at the
--         beginning of the processing stage, to allow for any hardware setup.
--
-- [start]: Signal which is asserted for as long as the processing stage is active.
--          Will remain high until [done] is asserted.
--
-- [btn_X]: These four signals are mapped to their corresponding buttons
--          on the FPGA development board. By default, left and right are
--          used by the transceiver to display the delay counter on the LEDs.
--          In order to utilize the LEDs for your hardware, you must assert
--          [override_leds] when a button is pressed and set [leds] as desired.
--
-- [switches]: The 16 dip switches on the FPGA development board.
--
-- [input]: Parallel input of size [G_total_bits] from the transceiver.
--
-- [output]: Parallel output of size [G_total_bits] back to the transceiver.
--
-- [done]: Done signal for the transceiver to terminate the processing stage
--         and begin to transmit the result (from [output]) back over UART.
--
-- [override_leds]: Signal to use [leds] from the hardware instead of transceiver.
--
-- [leds]: Output LEDs. Controlled by the top-level component based on [override_leds].
--
-------------------------------------------------------------------------------------

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
  use IEEE.std_logic_unsigned.all;
  use IEEE.math_real.all;

entity hw_container is
  generic (
    G_byte_bits  : integer := 8;
    G_total_bits : integer := 128;
    G_clk_freq   : integer := 100_000_000
  );
  port (
    clk_100mhz    : in    std_logic; -- board clk
    clk_hw        : in    std_logic; -- clock to be passed to hardware
    reset         : in    std_logic; -- async reset which is high when xcvr is not in processing stage
    load          : in    std_logic; -- pseudo-async pulse received from xcvr at the start of processing stage
    start         : in    std_logic; -- consistent signal received from xcvr as long as processing stage is active
    btn_up        : in    std_logic;
    btn_left      : in    std_logic; -- left is by default used for displaying left half of delay counter from xcvr
    btn_right     : in    std_logic; -- right is by default used for displaying right half of delay counter from xcvr
    btn_down      : in    std_logic;
    switches      : in    std_logic_vector(15 downto 0);
    input         : in    std_logic_vector(G_total_bits - 1 downto 0);
    output        : out   std_logic_vector(G_total_bits - 1 downto 0);
    done          : out   std_logic; -- tells xcvr to finish processing stage and transmit back result ([output])
    override_leds : out   std_logic; -- tells xcvr to use [leds] instead of displaying bytes received or delay
    leds          : out   std_logic_vector(15 downto 0)
  );
end hw_container;

architecture behavioral of hw_container is

  signal hw_done  : std_logic;
  signal leds_buf : std_logic_vector(15 downto 0);

  signal sum    : std_logic_vector(63 downto 0);
  signal c_out  : std_logic;

  signal s_mr   : std_logic;
  signal s_md   : std_logic;
  signal s_prod : std_logic;
  
  component cla_pow_4 is
    generic (
      G_size : integer
    );
    port (
      a      : in    std_logic_vector(G_size - 1 downto 0);
      b      : in    std_logic_vector(G_size - 1 downto 0);
      c_in   : in    std_logic;
      sum    : out   std_logic_vector(G_size - 1 downto 0);
      c_out  : out   std_logic;
      prop_g : out   std_logic;
      gen_g  : out   std_logic
    );
  end component;

  component two_level_multiplier is
    generic (
      G_n : integer := 64; -- Input (multiplier) length is n
      G_m : integer := 64  -- Input (multiplicand) length is m
    );
    port (
      clk    : in    std_logic;
      reset  : in    std_logic;
      start  : in    std_logic;
      s_mr   : in    std_logic;
      mr     : in    std_logic_vector(G_n - 1 downto 0);
      s_md   : in    std_logic;
      md     : in    std_logic_vector(G_m - 1 downto 0);
      s_prod : out   std_logic;
      prod   : out   std_logic_vector(G_n + G_m - 1 downto 0);
      done   : out   std_logic
    );
  end component;

  component d_flip_flop is
    port (
      input  : in    std_logic;
      clk    : in    std_logic;
      reset  : in    std_logic;
      output : out   std_logic
    );
  end component;

begin

  leds          <= leds_buf;
  done          <= hw_done;
  override_leds <= '1';

  ---------------------------------------------------------------------------
  -- Lab 12
  ---------------------------------------------------------------------------
  -- Uncomment the corresponding section of code during each part.
  -- Comment out the code for previous parts when advancing to the next.
  -- Tip: Select all lines in the section and press `CTRL + /` to do this.
  ---------------------------------------------------------------------------

  process (clk_hw, reset) begin
    if (reset = '1') then
      leds_buf <= (others => '0');
    elsif (clk_hw'event and clk_hw = '1') then
      if (start = '1' and hw_done = '0') then -- Only update while the hardware is running
        leds_buf(15)          <= s_prod;
        leds_buf(14 downto 2) <= (others => '0');
        leds_buf(1)           <= s_mr;
        leds_buf(0)           <= s_md;
      end if;
    end if;
  end process;

  --------------------------------------------
  -- Part B
  --------------------------------------------

--  adder : cla_pow_4
--    generic map (
--      G_size => 64
--    )
--    port map (
--      a      => input(127 downto 64),
--      b      => input(63 downto 0),
--      c_in   => '0',
--      sum    => sum,
--      c_out  => c_out,
--      prop_g => open,
--      gen_g  => open
--    );

--  done_generator : d_flip_flop
--    port map (
--      input  => start,
--      clk    => clk_hw,
--      reset  => reset,
--      output => hw_done
--    );
  
--  output(63 downto 0) <= sum; 
--  output(64) <= c_out;
--  output(output'left downto 65) <= (others => '0');

  --------------------------------------------
  -- Part C
  --------------------------------------------

   s_mr <= switches(1);
   s_md <= switches(0);

   multiplier : two_level_multiplier
     generic map (
       G_n => 64,
       G_m => 64
     )
     port map (
       clk    => clk_hw,
       reset  => reset,
       start  => start,
       s_mr   => s_mr,
       mr     => input(127 downto 64),
       s_md   => s_md,
       md     => input(63 downto 0),
       s_prod => s_prod,
       prod   => output,
       done   => hw_done
     );

end architecture behavioral;
