----------------------------------------------------------------------------
-- mk8_apex_128.vhd
----------------------------------------------------------------------------
-- Author:      Maxwell Phillips
-- Copyright:   Ohio Northern University, 2023.
-- License:     GPL v3
-- Description: Apex Component Linking Module
----------------------------------------------------------------------------
--
-- This file is a top-level component primarily designed for using a
-- serial UART RS-232 transceiver and an arbitrary hardware component,
-- such as a high-precision multiplier, alongside a Xilinx MMCM/PLL IP
-- core generated by the Vivado Clock Wizard. You will need to create
-- and customize the IP core appropriately for your design and link
-- its outputs to the appropriate ports and subcomponents.
--
----------------------------------------------------------------------------
-- Modification for Arbitrary Precisions
----------------------------------------------------------------------------
--
-- Change [G_total_bits] to desired precision.
-- It is recommended to change the filename as well (ex. mk8_apex_1024.vhd).
--
----------------------------------------------------------------------------
-- Modification for Arbitrary Hardware
----------------------------------------------------------------------------
--
-- Modify the `hw_container` component internally as appropriate.
-- You should not have to change this file for different hardwares, except
-- perhaps to increase the number of flip-flops for CDC synchronization.
-- To change hardware clock rate, re-customize the `hw_mmcm` (clk_wiz_0) IP.
--
----------------------------------------------------------------------------
-- Generics
----------------------------------------------------------------------------
--
-- [G_byte_bits]: Number of bits in a byte. Should be 8. Do not change.
--
-- [G_total_bits]: The capacity, in bits, of the transceiver and hardware.
--
-- [G_clk_freq]: Should match the clock frequency of the FPGA board (100 MHz).
--
-- [G_sampling_factor]: Factor to oversample by when receiving. Recommended 4-16.
--
-- [G_baud_rate]: Standard baud rate to use. Default 9600.
--
----------------------------------------------------------------------------
-- Ports
----------------------------------------------------------------------------
--
-- [clk]: Input clock signal; should match [G_clk_freq] generic.
--
-- [reset]: Asynchronous reset signal. This component also has an
--          initial reset signal built-in. This is mapped to the
--          center button on the FPGA development board.
--
-- [btn_X]: These four signals are mapped to their corresponding buttons
--          on the FPGA development board. They are passed to the transceiver
--          and the hardware container.
--
-- [switches]: The (16) dip switches on the FPGA development board.
--             Passed through to hardware container.
--
-- [input]: Serial UART input pin. Constrain appropriately. Passed to XCVR/RX.
--
-- [output]: Serial UART output pin. Constrain appropriately. Passed to XCVR/TX.
--
-- [leds]: The (16) LEDs on the FPGA development board.
--         Controlled by the transceiver and hardware container.
--
----------------------------------------------------------------------------

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
  use IEEE.std_logic_unsigned.all;

entity apex is
  generic (
    G_byte_bits       : integer := 8;           -- # of bits in a byte. do not change.
    G_total_bits      : integer := 128;        -- input length
    G_clk_freq        : integer := 100_000_000; -- board clk
    G_sampling_factor : integer := 4;           -- rx oversampling factor
    G_baud_rate       : integer := 9600
  );
  port (
    clk       : in    std_logic;
    reset     : in    std_logic;
    btn_up    : in    std_logic;
    btn_left  : in    std_logic;
    btn_right : in    std_logic;
    btn_down  : in    std_logic;
    switches  : in    std_logic_vector(15 downto 0);
    input     : in    std_logic; -- serial in
    output    : out   std_logic; -- serial out
    leds      : out   std_logic_vector(15 downto 0)
  );
end apex;

architecture behavioral of apex is

  --------------------------
  -- Clock Wizard IP Core --
  --------------------------

  component clk_wiz_0 is
    port (
      reset      : in    std_logic;
      clk_in1    : in    std_logic;
      clk_100mhz : out   std_logic;
      clk_hw     : out   std_logic;
      locked     : out   std_logic
    );
  end component;

  signal mmcm_locked : std_logic;
  signal clk_100mhz  : std_logic;
  signal clk_hw      : std_logic;
  signal clk_hw_buf  : std_logic;

  -----------------
  -- Transceiver --
  -----------------

  constant G_bytes : integer := G_total_bits / G_byte_bits;

  component transceiver is
    generic (
      G_byte_bits       : integer;
      G_bytes           : integer;
      G_total_bits      : integer;
      G_clk_freq        : integer;
      G_sampling_factor : integer;
      G_baud_rate       : integer
    );
    port (
      clk       : in    std_logic;
      reset     : in    std_logic;
      btn_up    : in    std_logic;
      btn_left  : in    std_logic;
      btn_right : in    std_logic;
      btn_down  : in    std_logic;
      switches  : in    std_logic_vector(15 downto 0);
      input     : in    std_logic;
      output    : out   std_logic;
      leds      : out   std_logic_vector(15 downto 0);

      -- HW Container Linkage
      data_out         : out   std_logic_vector(G_total_bits - 1 downto 0);
      hw_reset         : out   std_logic;
      hw_load          : out   std_logic;
      hw_start         : out   std_logic;
      hw_done          : in    std_logic;
      hw_output        : in    std_logic_vector(G_total_bits - 1 downto 0)
    );
  end component;

  signal xcvr_reset : std_logic;
  signal xcvr_data  : std_logic_vector(G_total_bits - 1 downto 0);
  signal xcvr_leds  : std_logic_vector(15 downto 0);

  ------------------------
  -- Hardware Container --
  ------------------------

  component hw_container is
    generic (
      G_byte_bits  : integer;
      G_clk_freq   : integer;
      G_total_bits : integer
    );
    port (
      clk_100mhz    : in    std_logic;
      clk_hw        : in    std_logic;
      reset         : in    std_logic;
      load          : in    std_logic;
      start         : in    std_logic;
      btn_up        : in    std_logic;
      btn_left      : in    std_logic;
      btn_right     : in    std_logic;
      btn_down      : in    std_logic;
      switches      : in    std_logic_vector(15 downto 0);
      input         : in    std_logic_vector(G_total_bits - 1 downto 0);
      output        : out   std_logic_vector(G_total_bits - 1 downto 0);
      done          : out   std_logic;
      override_leds : out   std_logic;
      leds          : out   std_logic_vector(15 downto 0)
    );
  end component;

  signal hw_reset         : std_logic;
  signal hw_load          : std_logic;
  signal hw_start         : std_logic;
  signal hw_start_sync    : std_logic;
  signal hw_done          : std_logic;
  signal hw_done_sync     : std_logic;
  signal hw_output        : std_logic_vector(G_total_bits - 1 downto 0);
  signal hw_leds          : std_logic_vector(15 downto 0);
  signal hw_override_leds : std_logic;

  component d_flip_flop is
    port (
      input  : in    std_logic;
      clk    : in    std_logic;
      reset  : in    std_logic;
      output : out   std_logic
    );
  end component;

  component synchronizer_2ff is
    port (
      input    : in    std_logic;
      dest_clk : in    std_logic;
      reset    : in    std_logic;
      output   : out   std_logic
    );
  end component; 

begin

  leds <= hw_leds when (hw_override_leds = '1') else xcvr_leds;

  xcvr_reset <= reset;

  hw_mmcm : clk_wiz_0
    port map (
      reset      => reset,
      clk_in1    => clk,
      clk_100mhz => clk_100mhz,
      clk_hw     => clk_hw_buf,
      locked     => mmcm_locked
    );

  clk_hw <= clk_hw_buf when (mmcm_locked = '1') else '0';

  xcvr : transceiver
    generic map (
      G_byte_bits       => G_byte_bits,
      G_bytes           => G_bytes,
      G_total_bits      => G_total_bits,
      G_clk_freq        => G_clk_freq,
      G_sampling_factor => G_sampling_factor,
      G_baud_rate       => G_baud_rate
    )
    port map (
      clk              => clk,
      reset            => xcvr_reset,
      btn_up           => btn_up,
      btn_left         => btn_left,
      btn_right        => btn_right,
      btn_down         => btn_down,
      switches         => switches,
      input            => input,
      output           => output,
      leds             => xcvr_leds,
      data_out         => xcvr_data,
      hw_reset         => hw_reset,
      hw_load          => hw_load,
      hw_start         => hw_start,
      hw_done          => hw_done_sync,
      hw_output        => hw_output
    );

  hw : hw_container
    generic map (
      G_byte_bits  => G_byte_bits,
      G_total_bits => G_total_bits,
      G_clk_freq   => G_clk_freq
    )
    port map (
      clk_100mhz    => clk,
      clk_hw        => clk_hw,
      reset         => hw_reset,
      load          => hw_load,
      start         => hw_start_sync,
      btn_up        => btn_up,
      btn_left      => btn_left,
      btn_right     => btn_right,
      btn_down      => btn_down,
      switches      => switches,
      input         => xcvr_data,
      output        => hw_output,
      done          => hw_done,
      override_leds => hw_override_leds,
      leds          => hw_leds
    );

  start_syncr : synchronizer_2ff
    port map (
      input    => hw_start,
      dest_clk => clk_hw,
      reset    => reset,
      output   => hw_start_sync
    );

  done_syncr : synchronizer_2ff
    port map (
      input    => hw_done,
      dest_clk => clk,
      reset    => reset,
      output   => hw_done_sync
    );

end architecture behavioral;
