-------------------------------------------------------------------------------------
-- Transceiver Hardware Component Container, version 2 (for Mk8 Apex/XCVR)
-------------------------------------------------------------------------------------
-- Author:      Maxwell Phillips
-- Copyright:   Ohio Northern University, 2023.
-- License:     GPL v3
-- Description: Container for hardware to be wrapped by apex component.
-------------------------------------------------------------------------------------
--
-- This file is the hardware component container wrapped by the top level apex 
-- component. You should modify this file to wrap your hardware in order to utilize
-- it with the serial transceiver. See the apex component and transceiver files
-- for more details on their functionality.
--
-------------------------------------------------------------------------------------
-- Generics
-------------------------------------------------------------------------------------
--
-- [G_byte_bits]: Should be 8. Mapped from top-level component.
--
-- [G_total_bits]: The capacity, in bits, of the transceiver. 
--                 Mapped directly from the top-level component.
--                 Should be used to help structure hardware components.
--
-- [G_clk_freq]: Should match the clock frequency of the FPGA board.
--               Again, mapped by top-level component.
--
-------------------------------------------------------------------------------------
-- Ports
-------------------------------------------------------------------------------------
--
-- [clk_100mhz]: Input clock signal; should match [G_clk_freq] generic.
--
-- [clk_hw]: Clock signal to time contained hardware. Generated by MMCM on top-level.
--
-- [reset]: Asynchronous reset signal. The module should be initially 
--          reset automatically by the transceiver, and will remain reset
--          until all bytes are received and the processing stage begins.
--          To preserve state, the hardware is NOT reset after the processing
--          stage and during the transmission stage. This allows displaying
--          output on the LEDs from the hardware container more easily.
--
-- [load]: Signal which is received for one clock cycle (of [G_clk_freq]) at the 
--         beginning of the processing stage, to allow for any hardware setup.
--
-- [start]: Signal which is asserted for as long as the processing stage is active.
--          Will remain high until [done] is asserted.
--
-- [btn_X]: These four signals are mapped to their corresponding buttons
--          on the FPGA development board. By default, left and right are 
--          used by the transceiver to display the delay counter on the LEDs.
--          In order to utilize the LEDs for your hardware, you must assert
--          [override_leds] when a button is pressed and set [leds] as desired. 
--
-- [switches]: The 16 dip switches on the FPGA development board. 
--
-- [input]: Parallel input of size [G_total_bits] from the transceiver.
-- 
-- [output]: Parallel output of size [G_total_bits] back to the transceiver.
--
-- [done]: Done signal for the transceiver to terminate the processing stage
--         and begin to transmit the result (from [output]) back over UART.
--
-- [override_leds]: Signal to use [leds] from the hardware instead of transceiver.
--
-- [leds]: Output LEDs. Controlled by the top-level component based on [override_leds].
--
-------------------------------------------------------------------------------------

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
  use IEEE.std_logic_unsigned.all;
  use IEEE.math_real.all;

entity hw_container is
  generic (
    G_byte_bits  : integer := 8;
    G_total_bits : integer := 64;
    G_clk_freq   : integer := 100_000_000
  );
  port (
    clk_100mhz    : in    std_logic; -- board clk
    clk_hw        : in    std_logic; -- clock to be passed to hardware
    reset         : in    std_logic; -- async reset which is high when xcvr is not in processing stage
    load          : in    std_logic; -- pseudo-async pulse received from xcvr at the start of processing stage
    start         : in    std_logic; -- consistent signal received from xcvr as long as processing stage is active
    btn_up        : in    std_logic;
    btn_left      : in    std_logic; -- left is by default used for displaying left half of delay counter from xcvr
    btn_right     : in    std_logic; -- right is by default used for displaying right half of delay counter from xcvr
    btn_down      : in    std_logic;
    switches      : in    std_logic_vector(15 downto 0);
    input         : in    std_logic_vector(G_total_bits - 1 downto 0);
    output        : out   std_logic_vector(G_total_bits - 1 downto 0);
    done          : out   std_logic; -- tells xcvr to finish processing stage and transmit back result ([output])
    override_leds : out   std_logic; -- tells xcvr to use [leds] instead of displaying bytes received or delay
    leds          : out   std_logic_vector(15 downto 0)
  );
end entity hw_container;

architecture behavioral of hw_container is

  constant G_n       : integer := G_total_bits;
  constant G_log_2_n : integer := integer(round(log2(real(G_n))));                  -- Base 2 Logarithm of input length n
  constant G_q       : integer := integer(round(2 ** ceil(log2(sqrt(real(G_n)))))); -- q is the least power of 2 greater than sqrt(n).
  constant G_log_2_q : integer := integer(round(log2(real(G_q))));                  -- Base 2 Logarithm of q
  constant G_k       : integer := G_n / G_q;                                        -- k is defined as n/q, if n is a perfect square, then k = sqrt(n) = q
  constant G_log_2_k : integer := integer(round(log2(real(G_k))));                  -- Base 2 Logarithm of k

  component priority_encoder_64 is
    port (
      input  : in    std_logic_vector(G_n - 1 downto 0);
      output : out   std_logic_vector(G_log_2_n - 1 downto 0);
      valid  : out   std_logic
    );
  end component priority_encoder_64;

  component barrel_shifter_generic is
    generic (
      G_n       : integer;
      G_log_2_n : integer;
      G_m       : integer;
      G_q       : integer;
      G_log_2_q : integer;
      G_k       : integer;
      G_log_2_k : integer
    );
    port (
      input  : in    std_logic_vector(G_n - 1 downto 0);
      shamt  : in    std_logic_vector(G_log_2_n - 1 downto 0);
      output : out   std_logic_vector(2 * G_n - 1 downto 0)
    );
  end component barrel_shifter_generic;

  component decoder_generic is
    generic (
      G_input_size  : integer;
      G_coarse_size : integer;
      G_fine_size   : integer
    );
    port (
      input  : in    std_logic_vector(G_input_size - 1 downto 0);
      output : out   std_logic_vector((2 ** G_input_size) - 1 downto 0)
    );
  end component decoder_generic;

  signal encoder_valid  : std_logic;
  signal encoder_output : std_logic_vector(G_log_2_n - 1 downto 0);
  signal shifter_output : std_logic_vector(2 * G_n - 1 downto 0);
  signal hw_done        : std_logic;
  signal leds_buf       : std_logic_vector(15 downto 0);
  signal dff1_out       : std_logic;

  component d_flip_flop is
    port (
      input  : in    std_logic;
      clk    : in    std_logic;
      reset  : in    std_logic;
      output : out   std_logic
    );
  end component;

begin

  done_generator : d_flip_flop
    port map (
      input  => start,
      clk    => clk_hw,
      reset  => reset,
      output => hw_done
    );

  leds <= leds_buf;
  done <= hw_done;
  override_leds <= '1';

  ---------------------------------------------------------------------------
  -- Lab 11                                                       
  ---------------------------------------------------------------------------
  -- Uncomment the corresponding section of code during each part.
  -- Comment out the code for previous parts when advancing to the next.
  -- Tip: Select all lines in the section and press `CTRL + /` to do this.
  ---------------------------------------------------------------------------

  process (clk_hw, reset) begin
    if (reset = '1') then
      leds_buf <= (others => '0');
    elsif (clk_hw'event and clk_hw = '1') then
        
        --------------------------------------------
        -- Part B, Section 1
        --------------------------------------------

        if (start = '1' and hw_done = '0') then -- Only update while the hardware is running
          leds_buf <= (15 => encoder_valid, others => '0');
        end if;        

        --------------------------------------------
        -- Part D, Section 1
        --------------------------------------------

        -- if (start = '1' and hw_done = '0') then -- Only update while the hardware is running
        --   leds_buf <= (G_log_2_n - 1 downto 0 => switches(G_log_2_n - 1 downto 0), others => '0');
        -- end if;
        
    end if;
  end process;
  
  --------------------------------------------
  -- Part B, Section 2
  --------------------------------------------

  encoder : priority_encoder_64
    port map (
      input  => input,
      output => encoder_output,
      valid  => encoder_valid
    );

  output <= (G_log_2_n - 1 downto 0 => encoder_output, others => '0');

  --------------------------------------------
  -- Part C
  --------------------------------------------

  -- decoder : decoder_generic
  --   generic map (
  --     G_input_size  => G_log_2_n,
  --     G_coarse_size => G_log_2_k,
  --     G_fine_size   => G_log_2_q
  --   )
  --   port map (
  --     input  => input(G_log_2_n - 1 downto 0),
  --     output => output
  --   );

  --------------------------------------------
  -- Part D, Section 2
  --------------------------------------------

  -- shifter : barrel_shifter_generic
  --   generic map (
  --     G_n       => G_n,
  --     G_log_2_n => G_log_2_n,
  --     G_m       => G_n,
  --     G_q       => G_q,
  --     G_log_2_q => G_log_2_q,
  --     G_k       => G_k,
  --     G_log_2_k => G_log_2_k
  --   )
  --   port map (
  --     input  => input,
  --     shamt  => switches(5 downto 0),
  --     output => shifter_output
  --   );

  -- output <= shifter_output(G_n - 1 downto 0);

end architecture behavioral;
